** Profile: "NMOS_TRANSIENT_ANALYSIS-transient_analysis"  [ C:\Users\Public\Downloads\CAD\MOSFET-PSpiceFiles\NMOS_TRANSIENT_ANALYSIS\transient_analysis.sim ] 

** Creating circuit file "transient_analysis.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Cadence\SPB_16.5\tools\PSpice\PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.TRAN  0 8us 0 
.PROBE V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\NMOS_TRANSIENT_ANALYSIS.net" 


.END
