** Profile: "INVERTER-input_characterstics"  [ C:\Users\Public\Downloads\CAD\MOSFET-PSpiceFiles\INVERTER\input_characterstics.sim ] 

** Creating circuit file "input_characterstics.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\Cadence\SPB_16.5\tools\PSpice\PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.DC LIN V_V2 0 10 0.005 
+ LIN V_V1 0 5 1 
.PROBE V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\INVERTER.net" 


.END
